module Ship_Sprites(
	input logic 	[9:0] DrawX, DrawY,
	output logic	[7:0] ShipR, ShipG, ShipB
);

parameter bit [7:0] SpriteTableR[18:0][16:0] = '{
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'hff,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'hff,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'hff,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'hff,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'hde,8'hde,8'hde,8'hde,8'hde,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'hff,8'h00,8'h00,8'hde,8'h00,8'hde,8'hde,8'hff,8'hde,8'hde,8'h00,8'hde,8'h00,8'h00,8'hff,8'h00},
'{8'h00,8'hff,8'h00,8'h00,8'h00,8'hde,8'hde,8'hff,8'hff,8'hff,8'hde,8'hde,8'h00,8'h00,8'h00,8'hff,8'h00},
'{8'h00,8'hde,8'h00,8'h00,8'hde,8'hde,8'hde,8'hff,8'hde,8'hff,8'hde,8'hde,8'hde,8'h00,8'h00,8'hde,8'h00},
'{8'h00,8'hde,8'h00,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h00,8'hde,8'h00},
'{8'h00,8'hde,8'hde,8'hde,8'hde,8'hde,8'hff,8'hde,8'hde,8'hde,8'hff,8'hde,8'hde,8'hde,8'hde,8'hde,8'h00},
'{8'h00,8'hde,8'hde,8'hde,8'h00,8'hff,8'hff,8'hde,8'hde,8'hde,8'hff,8'hff,8'h00,8'hde,8'hde,8'hde,8'h00},
'{8'h00,8'hde,8'hde,8'h00,8'h00,8'hff,8'hff,8'h00,8'hde,8'h00,8'hff,8'hff,8'h00,8'h00,8'hde,8'hde,8'h00},
'{8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}
};

parameter bit [7:0] SpriteTableG[18:0][16:0] = '{
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}, 
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}, 
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}, 
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}, 
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}, 
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}, 
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}, 
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}, 
'{8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'hde,8'hde,8'hde,8'hde,8'hde,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00}, 
'{8'h00,8'h00,8'h00,8'h00,8'hde,8'h68,8'hde,8'hde,8'h00,8'hde,8'hde,8'h68,8'hde,8'h00,8'h00,8'h00,8'h00}, 
'{8'h00,8'h00,8'h00,8'h00,8'h68,8'hde,8'hde,8'h00,8'h00,8'h00,8'hde,8'hde,8'h68,8'h00,8'h00,8'h00,8'h00}, 
'{8'h00,8'hde,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'hde,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'hde,8'h00}, 
'{8'h00,8'hde,8'h00,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h00,8'hde,8'h00}, 
'{8'h00,8'hde,8'hde,8'hde,8'hde,8'hde,8'h00,8'hde,8'hde,8'hde,8'h00,8'hde,8'hde,8'hde,8'hde,8'hde,8'h00}, 
'{8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00}, 
'{8'h00,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'h00}, 
'{8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00}, 
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}, 
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}
};

parameter bit [7:0] SpriteTableB[18:0][16:0] = '{
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00, 8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00, 8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00, 8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00, 8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00, 8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00, 8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00, 8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00, 8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'hde,8'hde,8'hde,8'hde,8'hde,8'h00,8'hde,8'h00,8'h00,8'h00, 8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'hde,8'h00,8'hde,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00, 8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'h00,8'h00,8'h00,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00, 8'h00},
'{8'h00,8'hde,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'hde,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'hde, 8'h00},
'{8'h00,8'hde,8'h00,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h00,8'hde, 8'h00},
'{8'h00,8'hde,8'hde,8'hde,8'hde,8'hde,8'h00,8'hde,8'hde,8'hde,8'h00,8'hde,8'hde,8'hde,8'hde,8'hde, 8'h00},
'{8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde, 8'h00},
'{8'h00,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde, 8'h00},
'{8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde, 8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00, 8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00, 8'h00}
};

assign ShipR = SpriteTableR[DrawY][DrawX];
assign ShipG = SpriteTableG[DrawY][DrawX];
assign ShipB = SpriteTableB[DrawY][DrawX];

endmodule

module Ship_Sprites2(
	input logic 	[9:0] DrawX, DrawY,
	output logic	[7:0] ShipR, ShipG, ShipB
);

parameter bit [7:0] SpriteTableR[18:0][16:0] = '{
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00, 8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00, 8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00, 8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00, 8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00, 8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00, 8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00, 8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00, 8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'hde,8'hde,8'hde,8'hde,8'hde,8'h00,8'hde,8'h00,8'h00,8'h00, 8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'hde,8'h00,8'hde,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00, 8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'h00,8'h00,8'h00,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00, 8'h00},
'{8'h00,8'hde,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'hde,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'hde, 8'h00},
'{8'h00,8'hde,8'h00,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h00,8'hde, 8'h00},
'{8'h00,8'hde,8'hde,8'hde,8'hde,8'hde,8'h00,8'hde,8'hde,8'hde,8'h00,8'hde,8'hde,8'hde,8'hde,8'hde, 8'h00},
'{8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde, 8'h00},
'{8'h00,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde, 8'h00},
'{8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde, 8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00, 8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00, 8'h00}
};

parameter bit [7:0] SpriteTableG[18:0][16:0] = '{
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}, 
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}, 
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}, 
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}, 
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}, 
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}, 
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}, 
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}, 
'{8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'hde,8'hde,8'hde,8'hde,8'hde,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00}, 
'{8'h00,8'h00,8'h00,8'h00,8'hde,8'h68,8'hde,8'hde,8'h00,8'hde,8'hde,8'h68,8'hde,8'h00,8'h00,8'h00,8'h00}, 
'{8'h00,8'h00,8'h00,8'h00,8'h68,8'hde,8'hde,8'h00,8'h00,8'h00,8'hde,8'hde,8'h68,8'h00,8'h00,8'h00,8'h00}, 
'{8'h00,8'hde,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'hde,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'hde,8'h00}, 
'{8'h00,8'hde,8'h00,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h00,8'hde,8'h00}, 
'{8'h00,8'hde,8'hde,8'hde,8'hde,8'hde,8'h00,8'hde,8'hde,8'hde,8'h00,8'hde,8'hde,8'hde,8'hde,8'hde,8'h00}, 
'{8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00}, 
'{8'h00,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'h00}, 
'{8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00}, 
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}, 
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}
};

parameter bit [7:0] SpriteTableB[18:0][16:0] = '{
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'hff,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'hff,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'hff,8'h00,8'h00,8'hde,8'hde,8'hde,8'h00,8'h00,8'hff,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'hde,8'hde,8'hde,8'hde,8'hde,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'hff,8'h00,8'h00,8'hde,8'h00,8'hde,8'hde,8'hff,8'hde,8'hde,8'h00,8'hde,8'h00,8'h00,8'hff,8'h00},
'{8'h00,8'hff,8'h00,8'h00,8'h00,8'hde,8'hde,8'hff,8'hff,8'hff,8'hde,8'hde,8'h00,8'h00,8'h00,8'hff,8'h00},
'{8'h00,8'hde,8'h00,8'h00,8'hde,8'hde,8'hde,8'hff,8'hde,8'hff,8'hde,8'hde,8'hde,8'h00,8'h00,8'hde,8'h00},
'{8'h00,8'hde,8'h00,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h00,8'hde,8'h00},
'{8'h00,8'hde,8'hde,8'hde,8'hde,8'hde,8'hff,8'hde,8'hde,8'hde,8'hff,8'hde,8'hde,8'hde,8'hde,8'hde,8'h00},
'{8'h00,8'hde,8'hde,8'hde,8'h00,8'hff,8'hff,8'hde,8'hde,8'hde,8'hff,8'hff,8'h00,8'hde,8'hde,8'hde,8'h00},
'{8'h00,8'hde,8'hde,8'h00,8'h00,8'hff,8'hff,8'h00,8'hde,8'h00,8'hff,8'hff,8'h00,8'h00,8'hde,8'hde,8'h00},
'{8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hde,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}
};



assign ShipR = SpriteTableR[DrawY][DrawX];
assign ShipG = SpriteTableG[DrawY][DrawX];
assign ShipB = SpriteTableB[DrawY][DrawX];

endmodule
		
module ship_rocket(
	input logic [9:0]		DrawX, DrawY,
	output logic [7:0]	SRockR, SRockG, SRockB
);

parameter bit [7:0] SpriteTableR[7:0][2:0] = '{
'{8'h00,8'hff,8'h00},
'{8'h00,8'hff,8'h00},
'{8'hff,8'hff,8'hff},
'{8'hff,8'h00,8'hff},
'{8'h00,8'hde,8'h00},
'{8'h00,8'hde,8'h00},
'{8'h00,8'hde,8'h00},
'{8'h00,8'hde,8'h00}
};

parameter bit [7:0] SpriteTableG[7:0][2:0] = '{
'{8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00},
'{8'h00,8'hff,8'h00},
'{8'h00,8'hde,8'h00},
'{8'h00,8'hde,8'h00},
'{8'h00,8'hde,8'h00},
'{8'h00,8'hde,8'h00}
};

parameter bit [7:0] SpriteTableB[7:0][2:0] = '{
'{8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00},
'{8'h00,8'hde,8'h00},
'{8'h00,8'hde,8'h00},
'{8'h00,8'hde,8'h00},
'{8'h00,8'hde,8'h00},
'{8'h00,8'hde,8'h00}
};



assign SRockR = SpriteTableR[DrawY][DrawX];
assign SRockG = SpriteTableG[DrawY][DrawX];
assign SRockB = SpriteTableB[DrawY][DrawX];

endmodule 

module ship_rocket2(
	input logic [9:0]		DrawX, DrawY,
	output logic [7:0]	SRockR, SRockG, SRockB
);

parameter bit [7:0] SpriteTableR[7:0][2:0] = '{
'{8'h00,8'hff,8'h00},
'{8'h00,8'hff,8'h00},
'{8'hff,8'hff,8'hff},
'{8'hff,8'h00,8'hff},
'{8'h00,8'hde,8'h00},
'{8'h00,8'hde,8'h00},
'{8'h00,8'hde,8'h00},
'{8'h00,8'hde,8'h00}
};

parameter bit [7:0] SpriteTableG[7:0][2:0] = '{
'{8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00},
'{8'h00,8'hff,8'h00},
'{8'h00,8'hde,8'h00},
'{8'h00,8'hde,8'h00},
'{8'h00,8'hde,8'h00},
'{8'h00,8'hde,8'h00}
};

parameter bit [7:0] SpriteTableB[7:0][2:0] = '{
'{8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00},
'{8'h00,8'hde,8'h00},
'{8'h00,8'hde,8'h00},
'{8'h00,8'hde,8'h00},
'{8'h00,8'hde,8'h00},
'{8'h00,8'hde,8'h00}
};



assign SRockR = SpriteTableR[DrawY][DrawX];
assign SRockG = SpriteTableG[DrawY][DrawX];
assign SRockB = SpriteTableB[DrawY][DrawX];

endmodule 